
module top(
  input a,
  input b,
  output f
);
  assign f = a ^ b;
   // Print some stuff as an example
endmodule


